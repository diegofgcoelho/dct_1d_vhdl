library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.numeric_std.all;

package mypack is
    --Class A AI type
    subtype classA is signed(7 downto 0);
    --AI type
    type AI is array (0 to 7) of classA;
    --Class B AI type
    type classB is array (0 to 3) of classA;
    --Class C AI type
    type classC is array (0 to 1) of classA;
    --Class D AI type
    type classD is array (0 to 3) of classA;
    --Class E AI type 
    type classE is array (0 to 1) of classA;
    
    component in_rom_memory is
       port(
          clk: in std_logic;
          addr: in std_logic_vector(9 downto 0);
          data0: out signed(7 downto 0);
          data1: out signed(7 downto 0);
          data2: out signed(7 downto 0);
          data3: out signed(7 downto 0);
          data4: out signed(7 downto 0);
          data5: out signed(7 downto 0);
          data6: out signed(7 downto 0);
          data7: out signed(7 downto 0)         
       );
    end component;

    component out_rom_memory is
       port(
          clk: in std_logic;
          addr: in std_logic_vector(9 downto 0);
          data0: out signed(7 downto 0);
          data1: out signed(7 downto 0);
          data2: out signed(7 downto 0);
          data3: out signed(7 downto 0);
          data4: out signed(7 downto 0);
          data5: out signed(7 downto 0);
          data6: out signed(7 downto 0);
          data7: out signed(7 downto 0)
       );
    end component;

end mypack;

package body mypack is

function c_log2 (x : positive) return natural is
    variable i : natural;
    begin
        i := 0;  
        while (2**i < x) and i < 31 loop
            i := i + 1;
        end loop;
        return i;
end function;

end package body;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity in_rom_memory is
port(
    clk: in std_logic;
    addr: in std_logic_vector(9 downto 0);
    data0: out signed(7 downto 0);
    data1: out signed(7 downto 0);
    data2: out signed(7 downto 0);
    data3: out signed(7 downto 0);
    data4: out signed(7 downto 0);
    data5: out signed(7 downto 0);
    data6: out signed(7 downto 0);
    data7: out signed(7 downto 0)
    );
end in_rom_memory;

architecture arc of in_rom_memory is
   constant ADDR_WIDTH: integer:=10;
   constant DATA_WIDTH: integer:=8;
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant ROM: rom_type:=(  
"00001001",
   "00001100",
   "11110101",
   "00001100",
   "00000100",
   "11110100",
   "11111001",
   "00000001",
   "00001110",
   "00001110",
   "11110110",
   "00001110",
   "00001110",
   "00000000",
   "00001001",
   "11110101",
   "11111110",
   "00001100",
   "00001001",
   "00001110",
   "00000101",
   "11110010",
   "00001010",
   "00001101",
   "00000101",
   "00001000",
   "00000111",
   "11111101",
   "00000101",
   "11110110",
   "00000110",
   "11110010",
   "11111001",
   "11110010",
   "11110100",
   "00001010",
   "00000110",
   "11111011",
   "00001110",
   "11110010",
   "11111110",
   "11111100",
   "00001000",
   "00001001",
   "11110111",
   "00000000",
   "11111110",
   "00000100",
   "00000110",
   "00001000",
   "11111001",
   "00000101",
   "00000101",
   "11110110",
   "11110101",
   "00000000",
   "00001110",
   "11111011",
   "00000011",
   "11111000",
   "00001000",
   "11111001",
   "00000000",
   "00000110",
   "00001100",
   "00001110",
   "00000001",
   "11110101",
   "11110101",
   "11111001",
   "00001010",
   "11111001",
   "00001001",
   "11111000",
   "00001101",
   "11111011",
   "11110111",
   "11111001",
   "00000011",
   "11111111",
   "11111100",
   "00001010",
   "00000011",
   "00000001",
   "00001101",
   "11111010",
   "00001000",
   "00001000",
   "11111100",
   "00000010",
   "11110011",
   "11110011",
   "00000001",
   "00001000",
   "00001101",
   "11110101",
   "00000010",
   "11111111",
   "11110001",
   "11111011",
   "11110110",
   "00001001",
   "11111010",
   "00000001",
   "11110110",
   "00000011",
   "11111001",
   "00000101",
   "00000110",
   "00000111",
   "11111111",
   "11110100",
   "11111000",
   "00001100",
   "11110110",
   "00001010",
   "00000001",
   "00001111",
   "11110011",
   "11111110",
   "11110100",
   "00001110",
   "11110001",
   "00001000",
   "00001010",
   "00001011",
   "11110100",
   "11111101",
   "11111001",
   "00001001",
   "11111110",
   "00001100",
   "11110110",
   "11111001",
   "11110101",
   "11110101",
   "00001011",
   "00000010",
   "00000001",
   "11110101",
   "00001011",
   "00000100",
   "11111100",
   "00000000",
   "00001100",
   "00001101",
   "00000000",
   "00000000",
   "11111011",
   "00001100",
   "11111100",
   "11110100",
   "00000010",
   "11110011",
   "11111000",
   "11111100",
   "00001010",
   "11110001",
   "11110010",
   "11110110",
   "00000100",
   "00000111",
   "00000100",
   "11111111",
   "00000001",
   "11111010",
   "00000111",
   "11110111",
   "00000110",
   "11110111",
   "11111100",
   "00000100",
   "00001000",
   "11110011",
   "00001101",
   "00001000",
   "00000000",
   "11111110",
   "11111110",
   "11111010",
   "00000000",
   "00000000",
   "00001010",
   "00001001",
   "00000100",
   "11111100",
   "00001001",
   "00000001",
   "11111100",
   "00001101",
   "00001011",
   "00000010",
   "00000100",
   "00000011",
   "11110111",
   "11111010",
   "11111111",
   "11111000",
   "00001010",
   "11110111",
   "11111000",
   "11110110",
   "11111000",
   "11111110",
   "11111010",
   "00001101",
   "11111110",
   "11110111",
   "00001100",
   "00001110",
   "11111110",
   "11110100",
   "11111001",
   "11111101",
   "00000011",
   "11111001",
   "00000011",
   "00000110",
   "11111000",
   "11110101",
   "11111010",
   "11111011",
   "11111110",
   "00000000",
   "11110100",
   "11111001",
   "00001001",
   "11110010",
   "00001101",
   "00000111",
   "00000000",
   "00000010",
   "11111000",
   "11111111",
   "00001110",
   "00000001",
   "00000001",
   "11111000",
   "00000000",
   "00000100",
   "00000101",
   "11111101",
   "11111100",
   "00001111",
   "11110010",
   "00001100",
   "00001100",
   "00001001",
   "11110100",
   "11111001",
   "11111011",
   "00000101",
   "11110101",
   "00000111",
   "11110100",
   "00000101",
   "00000000",
   "00001000",
   "00000110",
   "00001100",
   "00001100",
   "11111011",
   "00000110",
   "11110111",
   "11110010",
   "00000111",
   "00000000",
   "11111111",
   "00001100",
   "00000011",
   "00000100",
   "00001011",
   "00001001",
   "00000010",
   "11110110",
   "11111000",
   "00001100",
   "11110010",
   "00000000",
   "11110110",
   "00001110",
   "00000110",
   "00000000",
   "11111111",
   "11110011",
   "00000101",
   "11110010",
   "11110011",
   "00000001",
   "11110100",
   "00001010",
   "00001010",
   "00000111",
   "11110101",
   "00000101",
   "00000001",
   "00001110",
   "00000100",
   "00001001",
   "11111111",
   "11111110",
   "00001010",
   "11110100",
   "11110101",
   "11110110",
   "11111101",
   "00001010",
   "00001001",
   "11110011",
   "11111101",
   "00000001",
   "11111110",
   "00000101",
   "00000100",
   "11111010",
   "11111110",
   "11110001",
   "00001111",
   "11110110",
   "11110100",
   "11111100",
   "11110111",
   "00000000",
   "11111011",
   "00001110",
   "00001101",
   "11110011",
   "00000111",
   "11111001",
   "11111110",
   "00000001",
   "00001101",
   "11111110",
   "00001110",
   "11111010",
   "00000110",
   "00000101",
   "00000001",
   "00000110",
   "00000101",
   "11110110",
   "11110101",
   "00001111",
   "11110110",
   "11110110",
   "00001011",
   "00000100",
   "11111100",
   "11110111",
   "11111110",
   "11111111",
   "11110101",
   "00000011",
   "11111000",
   "11111101",
   "00000010",
   "11111001",
   "11111010",
   "00000100",
   "11111001",
   "00001010",
   "00001110",
   "00000111",
   "11111011",
   "00000011",
   "11110100",
   "00001100",
   "00001011",
   "00001010",
   "11111001",
   "00000011",
   "11110010",
   "11111110",
   "11111010",
   "11110110",
   "11110110",
   "11111110",
   "11110100",
   "00000011",
   "11111111",
   "00000110",
   "00000110",
   "00000100",
   "11110010",
   "11110011",
   "11111011",
   "00000001",
   "00000101",
   "11111101",
   "00001010",
   "00000111",
   "00001110",
   "00000001",
   "11111011",
   "11110100",
   "00000011",
   "00001000",
   "11111110",
   "11110100",
   "11111001",
   "11110110",
   "11111001",
   "11111110",
   "00000001",
   "11111111",
   "00001011",
   "00000001",
   "00001101",
   "00000100",
   "00001110",
   "11111000",
   "00000101",
   "11111010",
   "00000101",
   "00000110",
   "11110011",
   "11111001",
   "11111000",
   "00000101",
   "00001010",
   "11111011",
   "00001000",
   "00000101",
   "11110001",
   "00000011",
   "11111101",
   "00001100",
   "11110001",
   "11111111",
   "11111110",
   "11111111",
   "00001000",
   "11111011",
   "00001001",
   "11111111",
   "11110010",
   "11110110",
   "00000111",
   "11111111",
   "11110110",
   "11111011",
   "00000011",
   "11110111",
   "00000111",
   "11111000",
   "00001101",
   "11111001",
   "00001000",
   "11110111",
   "11111010",
   "11110100",
   "00000010",
   "00000110",
   "00000001",
   "11111110",
   "00000100",
   "00000100",
   "00000101",
   "00000100",
   "00001101",
   "11110111",
   "00000110",
   "11111000",
   "11110101",
   "00000011",
   "11111111",
   "11111111",
   "00000101",
   "00001000",
   "11111100",
   "00000101",
   "11111101",
   "00001010",
   "00001010",
   "11111001",
   "00000011",
   "00000010",
   "00000001",
   "00001011",
   "11111001",
   "11111011",
   "11110101",
   "00001101",
   "00000100",
   "11111111",
   "00000100",
   "00000001",
   "00000100",
   "00000001",
   "00000111",
   "00000001",
   "00001111",
   "11111000",
   "11110100",
   "11110100",
   "11110011",
   "11111101",
   "11111110",
   "11111100",
   "00001000",
   "00000100",
   "00001000",
   "00001101",
   "00001110",
   "11110111",
   "11110101",
   "00000110",
   "11110100",
   "00000001",
   "00000001",
   "00001011",
   "00000000",
   "11111101",
   "00000101",
   "00000111",
   "00000001",
   "11111011",
   "11110101",
   "00000011",
   "11111001",
   "11110010",
   "00001000",
   "11111000",
   "11111110",
   "00000110",
   "11111100",
   "00000111",
   "11111101",
   "00000110",
   "00000110",
   "11111110",
   "11110010",
   "11111011",
   "11111110",
   "11111001",
   "11110111",
   "00001010",
   "11111110",
   "00001100",
   "11111101",
   "00001000",
   "11111101",
   "00001001",
   "00001000",
   "11111100",
   "11110111",
   "00001001",
   "00001101",
   "11111011",
   "00000101",
   "11111110",
   "00001010",
   "00001000",
   "11110110",
   "00001011",
   "00001111",
   "00000000",
   "00001100",
   "00000011",
   "11110110",
   "11110111",
   "11111101",
   "00000111",
   "00001010",
   "00001001",
   "11111011",
   "00000001",
   "11110100",
   "11110100",
   "11110101",
   "00000101",
   "00000000",
   "11110111",
   "00000000",
   "11110101",
   "11110011",
   "11110001",
   "00001011",
   "00000011",
   "00001111",
   "00000001",
   "11111111",
   "00001001",
   "11111000",
   "00000000",
   "00001100",
   "00000010",
   "00001010",
   "00000111",
   "00000011",
   "11111000",
   "00000101",
   "11110100",
   "00000100",
   "00000101",
   "00000111",
   "00001100",
   "00001110",
   "00001000",
   "00000010",
   "00000010",
   "00000100",
   "11110010",
   "00000011",
   "11111100",
   "11110010",
   "00000000",
   "11110111",
   "11110101",
   "11110111",
   "11110101",
   "11110111",
   "11110010",
   "00000100",
   "11111001",
   "00000001",
   "00000110",
   "00000000",
   "00000001",
   "11111110",
   "11110101",
   "00000000",
   "00001011",
   "00001011",
   "11111001",
   "11110111",
   "00000010",
   "00000100",
   "11111110",
   "11110111",
   "00001101",
   "11110011",
   "11110100",
   "11110101",
   "11110110",
   "00000100",
   "00000010",
   "11110011",
   "00001101",
   "00000111",
   "00000111",
   "11110011",
   "00001011",
   "00001101",
   "00001111",
   "00001011",
   "00001001",
   "00000000",
   "11110110",
   "11111101",
   "11110101",
   "11110010",
   "00001101",
   "11111010",
   "11111010",
   "11111011",
   "11111111",
   "00000100",
   "11110010",
   "00001010",
   "00000010",
   "00001011",
   "11111011",
   "11111110",
   "11110011",
   "11110110",
   "00000101",
   "11111011",
   "00001100",
   "11110101",
   "00001111",
   "00000001",
   "00000110",
   "00001111",
   "11111010",
   "11111101",
   "11111111",
   "00001000",
   "00001010",
   "11110100",
   "11110110",
   "11111100",
   "11110011",
   "00000001",
   "11111011",
   "11110110",
   "11110111",
   "00001100",
   "00000101",
   "11111111",
   "00001100",
   "11110100",
   "00000111",
   "00000111",
   "00000010",
   "11110111",
   "00000011",
   "11111010",
   "11110101",
   "11110111",
   "00001100",
   "11110011",
   "11111000",
   "11110011",
   "11111110",
   "11110001",
   "00001100",
   "11110111",
   "11110100",
   "11111010",
   "11111111",
   "11110100",
   "00001111",
   "11111011",
   "11111010",
   "11110011",
   "11111010",
   "11110010",
   "00000000",
   "00001000",
   "11111011",
   "11111010",
   "00000111",
   "11110001",
   "11110010",
   "00000101",
   "00000011",
   "00000001",
   "00000111",
   "00000110",
   "00001000",
   "11111010",
   "00000110",
   "00000010",
   "11111101",
   "11110011",
   "00001000",
   "11111011",
   "00000011",
   "00000111",
   "11110100",
   "11110101",
   "00000001",
   "00000000",
   "00000110",
   "11110101",
   "00000111",
   "11110100",
   "11110101",
   "00000100",
   "11111011",
   "00000101",
   "00000111",
   "00000010",
   "00000111",
   "11111000",
   "00000111",
   "00001110",
   "00001011",
   "11110100",
   "11111100",
   "11111100",
   "00000110",
   "00000011",
   "00001001",
   "11111100",
   "11110111",
   "11110100",
   "00001000",
   "11110111",
   "11111101",
   "00000010",
   "11111000",
   "00000100",
   "00000000",
   "11110110",
   "00001000",
   "11110100",
   "11111010",
   "11111000",
   "00000001",
   "11110100",
   "11111101",
   "11110100",
   "11110100",
   "00001001",
   "11111010",
   "00000011",
   "00001110",
   "11111110",
   "00000110",
   "00001000",
   "11111110",
   "00000101",
   "11110100",
   "00001101",
   "11110111",
   "11111001",
   "00001001",
   "00000000",
   "00001000",
   "11111101",
   "11111001",
   "11110010",
   "00000101",
   "11111110",
   "11111111",
   "00000011",
   "11110011",
   "11111010",
   "00001000",
   "00000110",
   "11110101",
   "11110101",
   "11110100",
   "11110001",
   "11111110",
   "00000101",
   "00000111",
   "00000001",
   "11110100",
   "00000100",
   "11110101",
   "11110101",
   "00001100",
   "00000110",
   "00000010",
   "11110111",
   "11110111",
   "11110011",
   "00001100",
   "00000110",
   "00000010",
   "11111010",
   "11110110",
   "00000100",
   "00001111",
   "11110110",
   "11111001",
   "11111101",
   "11110011",
   "00000110",
   "11111101",
   "00001110",
   "11111101",
   "00000100",
   "11110110",
   "11111100",
   "11110110",
   "00001000",
   "00001011",
   "11111100",
   "00000110",
   "11111010",
   "00000001",
   "00001010",
   "00000011",
   "11111011",
   "11111010",
   "11111111",
   "11111110",
   "11111100",
   "00000010",
   "00000111",
   "11111110",
   "11111110",
   "11110101",
   "11110010",
   "11111010",
   "11111011",
   "00000101",
   "00001110",
   "00001101",
   "11111111",
   "11111000",
   "00001000",
   "00001000",
   "00000111",
   "00000111",
   "11110100",
   "00000101",
   "11111111",
   "11110111",
   "11110100",
   "00001010",
   "11110110",
   "11110110",
   "00000101",
   "00001100",
   "00000000",
   "00000110",
   "11110110",
   "00001110",
   "00000001",
   "00000101",
   "11110010",
   "00001001",
   "00000111",
   "11110101",
   "00000001",
   "11111011",
   "00000001",
   "11111101",
   "11111101",
   "11110110",
   "11111001",
   "11110010",
   "00001101",
   "00000101",
   "00001101",
   "11110110",
   "00001101",
   "00001001",
   "00000010",
   "11111110",
   "11111001",
   "00001000",
   "11111000",
   "11110011",
   "00001000",
   "00000101",
   "00000110",
   "00000100",
   "11111110",
   "11111101",
   "00001001",
   "11111011",
   "00001001",
   "00001001",
   "00001011",
   "00000000",
   "00000100",
   "00001110",
   "11111110",
   "11110011",
   "00001011",
   "00000100",
   "11111100",
   "00001111",
   "11111000",
   "00000101",
   "00000011",
   "11111101",
   "11110101",
   "11110010",
   "11111110",
   "11110111",
   "00000111",
   "11111100",
   "00001010",
   "00000111",
   "00000010",
   "11110110",
   "00001110",
   "11111001",
   "00001101",
   "11111000",
   "11111100",
   "11110100",
   "00000100",
   "11110110",
   "11110010",
   "00000111",
   "11111011",
   "00000101",
   "11111101",
   "00000100",
   "11110010",
   "00001100",
   "00001001",
   "00000111",
   "00001001",
   "11111100",
   "00000100",
   "00000010",
   "00000001",
   "11111001",
   "11111000",
   "11111111",
   "11111000",
   "00001001",
   "00001111",
   "11110010",
   "00000001",
   "11110100",
   "00001001",
   "00001111",
   "11110011",
   "00001101",
   "11110010",
   "00000110",
   "00001001",
   "11110100",
   "00000011",
   "00001101",
   "11111100",
   "11111101",
   "00001111",
   "00001101",
   "00000101",
   "00001111",
   "00001000",
   "11111011",
   "00000101",
   "11111000",
   "11111010",
   "00000101",
   "00000001",
   "11111101",
   "00000011",
   "00001000",
   "00000011",
   "00000010",
   "00000011",
   "00000000",
   "11110011",
   "00000111",
   "00001111",
   "11111100",
   "00001110",
   "11111011",
   "00001100",
   "11111111",
   "11111101",
    others => "00000000"
   );
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (rising_edge(clk)) then
        addr_reg <= addr;
      end if;
   end process;
   data0 <= signed(ROM(to_integer(unsigned(addr_reg))));
   data1 <= signed(ROM(to_integer(unsigned(addr_reg))+1));
   data2 <= signed(ROM(to_integer(unsigned(addr_reg))+2));
   data3 <= signed(ROM(to_integer(unsigned(addr_reg))+3));
   data4 <= signed(ROM(to_integer(unsigned(addr_reg))+4));
   data5 <= signed(ROM(to_integer(unsigned(addr_reg))+5));
   data6 <= signed(ROM(to_integer(unsigned(addr_reg))+6));
   data7 <= signed(ROM(to_integer(unsigned(addr_reg))+7));
   
end arc;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity out_rom_memory is
port(
    clk: in std_logic;
    addr: in std_logic_vector(9 downto 0);
    data0: out signed(7 downto 0);
    data1: out signed(7 downto 0);
    data2: out signed(7 downto 0);
    data3: out signed(7 downto 0);
    data4: out signed(7 downto 0);
    data5: out signed(7 downto 0);
    data6: out signed(7 downto 0);
    data7: out signed(7 downto 0)

    );
end out_rom_memory;

architecture arc of out_rom_memory is
   constant ADDR_WIDTH: integer:=10;
   constant DATA_WIDTH: integer:=8;
   signal addr_reg: std_logic_vector(ADDR_WIDTH-1 downto 0);
   type rom_type is array (0 to 2**ADDR_WIDTH-1)
        of std_logic_vector(DATA_WIDTH-1 downto 0);
   -- ROM definition
   constant ROM: rom_type:=(  
"00010000",
   "01001000",
   "00001110",
   "11111000",
   "01011000",
   "11101011",
   "10110000",
   "11010010",
   "01011000",
   "01000001",
   "11100010",
   "01010011",
   "00100100",
   "00010011",
   "10001110",
   "11101110",
   "01011110",
   "00000100",
   "00001000",
   "10001101",
   "00011010",
   "00000100",
   "10110000",
   "00010001",
   "00001000",
   "01001111",
   "11110101",
   "00001000",
   "11011100",
   "00001110",
   "11000111",
   "01000101",
   "11010100",
   "11001000",
   "10110001",
   "00101101",
   "00011000",
   "01011110",
   "10101011",
   "00010100",
   "00001000",
   "00000001",
   "11110110",
   "11000000",
   "00000000",
   "00101010",
   "00100110",
   "11100000",
   "11111000",
   "01000010",
   "00000100",
   "11111011",
   "01001000",
   "11010110",
   "11010111",
   "11101100",
   "00010110",
   "00010001",
   "00110011",
   "00010010",
   "00111010",
   "11111010",
   "00011000",
   "01010000",
   "00000010",
   "01001010",
   "01100111",
   "00010100",
   "10111010",
   "00010111",
   "11001110",
   "00010111",
   "11110110",
   "00100011",
   "00101101",
   "11011111",
   "11110010",
   "01000010",
   "00110100",
   "00111010",
   "01000010",
   "11101010",
   "11111100",
   "11011100",
   "00000110",
   "11010000",
   "10111110",
   "00101100",
   "11011110",
   "11010000",
   "00001101",
   "01100110",
   "10110110",
   "11111101",
   "11001000",
   "00001010",
   "11001110",
   "11101011",
   "00101101",
   "00111010",
   "00000010",
   "11110010",
   "00010110",
   "10110010",
   "11101110",
   "11111000",
   "10101011",
   "00101010",
   "11100110",
   "11101101",
   "11010111",
   "11011100",
   "00001010",
   "00000111",
   "11000010",
   "00011011",
   "11111010",
   "10111000",
   "11111000",
   "10000001",
   "00000010",
   "11111010",
   "10110000",
   "00100111",
   "00001010",
   "10010110",
   "11001100",
   "10011010",
   "11001010",
   "01001110",
   "11010011",
   "11001101",
   "11110110",
   "00000101",
   "11011000",
   "10110001",
   "00011100",
   "00011011",
   "00010101",
   "01000001",
   "00010000",
   "11001011",
   "00011110",
   "00110010",
   "00100000",
   "01011010",
   "00001001",
   "01001000",
   "11001100",
   "11111011",
   "00001101",
   "11001000",
   "10011000",
   "00100110",
   "11010111",
   "00011110",
   "01100000",
   "11110011",
   "11111011",
   "00111100",
   "00001110",
   "00110010",
   "00000100",
   "00000101",
   "11011110",
   "00010101",
   "11010000",
   "00100100",
   "00011010",
   "11010010",
   "00011011",
   "11110100",
   "01001110",
   "00110101",
   "11001011",
   "01000001",
   "00010010",
   "11000100",
   "00110010",
   "00000000",
   "11111010",
   "00000011",
   "11110110",
   "00011001",
   "01000000",
   "11011110",
   "00000111",
   "00010000",
   "11001100",
   "00110110",
   "00110000",
   "00000001",
   "11100000",
   "00001111",
   "00100101",
   "00101101",
   "11110000",
   "00011011",
   "10110011",
   "00011101",
   "11000000",
   "11010001",
   "11010110",
   "00111010",
   "11011100",
   "00010101",
   "00100010",
   "11010000",
   "11111100",
   "01001101",
   "01010110",
   "00101011",
   "11001100",
   "11110100",
   "11100000",
   "00001001",
   "11010010",
   "00010011",
   "01000110",
   "00010010",
   "11110110",
   "11100001",
   "11101001",
   "11111011",
   "11111100",
   "10111100",
   "11001111",
   "00000111",
   "11011000",
   "10111111",
   "00110010",
   "01010010",
   "00000110",
   "11111110",
   "11101000",
   "10100111",
   "11110010",
   "11111100",
   "00001011",
   "00101110",
   "01000000",
   "11001000",
   "00100011",
   "11111101",
   "11111100",
   "01011110",
   "00001011",
   "10011111",
   "11000100",
   "11010010",
   "11100110",
   "11011101",
   "00001000",
   "11110110",
   "00110101",
   "10100110",
   "00111100",
   "00101110",
   "10110111",
   "11110101",
   "00000000",
   "00001110",
   "10111010",
   "00011011",
   "00101100",
   "10110101",
   "11100100",
   "11100000",
   "11110100",
   "10110000",
   "11011011",
   "00001010",
   "11011010",
   "00110100",
   "00001111",
   "00111111",
   "00110010",
   "11101011",
   "10110110",
   "01001000",
   "11100000",
   "01111000",
   "00011001",
   "00101111",
   "11101100",
   "00001100",
   "00110010",
   "11000010",
   "00010110",
   "11111010",
   "11010010",
   "11001010",
   "00110110",
   "01000001",
   "11111111",
   "01000011",
   "00010110",
   "01101001",
   "11110010",
   "00110011",
   "11101010",
   "11111100",
   "01001101",
   "11101111",
   "11101010",
   "00000000",
   "11100001",
   "10101000",
   "11010110",
   "00111001",
   "00001110",
   "11100011",
   "11010110",
   "00110110",
   "00001001",
   "01000110",
   "11001010",
   "00000110",
   "00110010",
   "10011101",
   "00000110",
   "11001011",
   "11001010",
   "00100101",
   "00101010",
   "10101111",
   "01010100",
   "00001001",
   "00100010",
   "11011001",
   "11000111",
   "11101011",
   "00000110",
   "11111100",
   "00101111",
   "10101010",
   "00000010",
   "00101011",
   "00010110",
   "11100100",
   "11010110",
   "01101011",
   "11001001",
   "00011100",
   "11010100",
   "00101011",
   "11110011",
   "11100011",
   "10100100",
   "11101111",
   "11100010",
   "11101101",
   "11010100",
   "00001001",
   "00001000",
   "00000111",
   "00001000",
   "01000111",
   "11110100",
   "00000110",
   "01010000",
   "00011011",
   "01011101",
   "11010100",
   "11111100",
   "11110000",
   "11000111",
   "00111111",
   "10111000",
   "01000110",
   "00011010",
   "00100111",
   "00001000",
   "11111111",
   "00110101",
   "00111100",
   "11101100",
   "11110011",
   "10110110",
   "00111000",
   "11101000",
   "00101101",
   "00010101",
   "00101100",
   "00100000",
   "10001111",
   "11110011",
   "11010011",
   "11101100",
   "00000100",
   "00010110",
   "11011000",
   "11001100",
   "00010100",
   "11010000",
   "00110010",
   "01001000",
   "11100111",
   "11110101",
   "11101111",
   "00001100",
   "10011010",
   "11110111",
   "11101111",
   "00000000",
   "11101111",
   "00101010",
   "11011011",
   "00001110",
   "00110011",
   "00000011",
   "00110110",
   "11001010",
   "00010111",
   "10111011",
   "10111111",
   "11110010",
   "11111011",
   "10101000",
   "00001010",
   "11001010",
   "01010010",
   "00001100",
   "11101000",
   "00000010",
   "11111011",
   "00110111",
   "11100100",
   "11101010",
   "11100100",
   "01000001",
   "01001000",
   "11001110",
   "00010110",
   "00011001",
   "00100010",
   "10010110",
   "11011110",
   "00000100",
   "11101011",
   "00000100",
   "11011001",
   "00000001",
   "00000001",
   "00000100",
   "11100110",
   "00011001",
   "10001011",
   "11100000",
   "10111011",
   "11100001",
   "00001101",
   "00101100",
   "11100110",
   "11101010",
   "11101011",
   "00001000",
   "01010001",
   "11010101",
   "11111111",
   "11101100",
   "00100110",
   "00010110",
   "10110010",
   "00011000",
   "00000101",
   "11100111",
   "00001101",
   "00011100",
   "00010100",
   "11011010",
   "00011100",
   "00101110",
   "00100000",
   "00011000",
   "00111101",
   "11110010",
   "00011011",
   "10110111",
   "11110101",
   "00010010",
   "11011011",
   "11011000",
   "11010000",
   "11110110",
   "00100011",
   "01000010",
   "00010101",
   "11010110",
   "01110100",
   "11010100",
   "11001110",
   "00010110",
   "00011110",
   "11011011",
   "11001000",
   "01001100",
   "10011100",
   "00000100",
   "11111011",
   "00010000",
   "00010001",
   "11101100",
   "11100110",
   "11100110",
   "10110011",
   "11111101",
   "11111101",
   "11001010",
   "00010011",
   "00010100",
   "01001101",
   "11101100",
   "00101111",
   "11111101",
   "11001100",
   "11011100",
   "00011000",
   "11011010",
   "00011000",
   "11101100",
   "11011001",
   "11100110",
   "11111101",
   "11100000",
   "11010110",
   "10100010",
   "00000101",
   "11001010",
   "01000011",
   "00101101",
   "00101010",
   "11011110",
   "11011110",
   "00001001",
   "00001100",
   "01001110",
   "11111101",
   "00011111",
   "11110010",
   "00001110",
   "00010000",
   "00010011",
   "01010100",
   "00100010",
   "11011000",
   "11011111",
   "10111011",
   "00010110",
   "00101001",
   "00111111",
   "11011010",
   "00111010",
   "00011010",
   "10110011",
   "00011100",
   "11111010",
   "01100011",
   "00111011",
   "11110010",
   "11111100",
   "00010010",
   "10010011",
   "11100110",
   "11111100",
   "00011000",
   "11011111",
   "00100001",
   "10011010",
   "00001111",
   "10111000",
   "11100110",
   "11011110",
   "00011001",
   "00110101",
   "11110011",
   "00011110",
   "11111111",
   "10101101",
   "11001101",
   "11000110",
   "00010010",
   "10100110",
   "11011011",
   "00111110",
   "00100001",
   "11011111",
   "11100111",
   "00011010",
   "11000111",
   "11110101",
   "11010011",
   "01010000",
   "10111110",
   "10101100",
   "00000010",
   "11010100",
   "11100100",
   "11110010",
   "11110111",
   "11000000",
   "00101011",
   "00010010",
   "00001100",
   "00100000",
   "00010110",
   "10100101",
   "11101100",
   "10010000",
   "11000101",
   "00011000",
   "00000110",
   "11101100",
   "11110110",
   "00100101",
   "11001011",
   "00100000",
   "11011110",
   "01011001",
   "11101001",
   "11110000",
   "00101100",
   "00000110",
   "11110111",
   "11010110",
   "11110001",
   "11010010",
   "11110010",
   "11100010",
   "01011010",
   "11001011",
   "00101111",
   "11011000",
   "10011000",
   "11111110",
   "11010101",
   "00101100",
   "00101011",
   "10110010",
   "00011100",
   "01101010",
   "11011110",
   "10101100",
   "00011111",
   "00100010",
   "01000011",
   "00101101",
   "00101011",
   "10101100",
   "11100010",
   "11100100",
   "00101010",
   "00010100",
   "10101101",
   "11011011",
   "00110111",
   "00001010",
   "11110101",
   "11011010",
   "00110110",
   "00011010",
   "11101101",
   "11101010",
   "10100001",
   "11110100",
   "10101110",
   "11011010",
   "11011011",
   "11111000",
   "00010000",
   "11001110",
   "01110100",
   "00100010",
   "00100110",
   "00010011",
   "01010001",
   "10110110",
   "00000001",
   "11000001",
   "11100110",
   "10110100",
   "11001101",
   "00011010",
   "11001000",
   "01000100",
   "11011100",
   "11101100",
   "11010100",
   "00010110",
   "00011101",
   "11101111",
   "00110010",
   "11000110",
   "11110100",
   "00110000",
   "01001100",
   "10100110",
   "00101000",
   "11101000",
   "00111111",
   "00111110",
   "11100011",
   "11010111",
   "01000100",
   "10100110",
   "00011000",
   "11111010",
   "11101000",
   "11001110",
   "01000111",
   "01000001",
   "00111101",
   "11010110",
   "00010000",
   "01111101",
   "00001000",
   "00111010",
   "00001100",
   "00000110",
   "00110001",
   "11010000",
   "11011100",
   "00110001",
   "11110010",
   "10101100",
   "00001110",
   "01000010",
   "00010010",
   "00001110",
   "01001111",
   "11101000",
   "00101100",
   "11011010",
   "11101101",
   "00001011",
   "00101100",
   "11101110",
   "00101000",
   "00100110",
   "11010001",
   "00011110",
   "01010001",
   "00000011",
   "11111010",
   "11011110",
   "11111000",
   "00111011",
   "11111110",
   "11110010",
   "00010001",
   "01101011",
   "00010011",
   "00111000",
   "00001100",
   "11101100",
   "01011100",
   "10110000",
   "00001111",
   "00010000",
   "00110001",
   "11100010",
   "00101110",
   "10100110",
   "11111101",
   "00001110",
   "11110110",
   "00001000",
   "00100100",
   "11100000",
   "00010111",
   "11111111",
   "00110011",
   "00000000",
   "01001000",
   "00011110",
   "11101011",
   "10101000",
   "00100110",
   "00001011",
   "00110001",
   "00101100",
   "00100110",
   "11111011",
   "01000000",
   "00101000",
   "11000011",
   "11100010",
   "11101011",
   "00001100",
   "10111100",
   "10101101",
   "00000101",
   "11111010",
   "11110101",
   "00010100",
   "11101000",
   "00001110",
   "00111000",
   "10100011",
   "10111100",
   "11101010",
   "11110110",
   "00111001",
   "00111000",
   "00011110",
   "11011101",
   "00001000",
   "00101110",
   "10010100",
   "00111010",
   "10110011",
   "10110001",
   "11101000",
   "00100100",
   "00001110",
   "11110101",
   "11011010",
   "01001010",
   "11101000",
   "11101111",
   "11000110",
   "00000001",
   "00101010",
   "11001110",
   "00001110",
   "00011010",
   "01111101",
   "11100111",
   "11110010",
   "00100010",
   "11011011",
   "00110000",
   "11100010",
   "00001010",
   "11010011",
   "00011100",
   "01100110",
   "11101011",
   "11011000",
   "00011111",
   "11101110",
   "00001011",
   "10110001",
   "11011010",
   "11111010",
   "11101001",
   "11101110",
   "10100010",
   "00100000",
   "11101110",
   "11111111",
   "10101101",
   "11101000",
   "10111111",
   "11110011",
   "00101101",
   "11110100",
   "11100001",
   "00101001",
   "11111110",
   "00101000",
   "00001110",
   "11111011",
   "00000001",
   "11010110",
   "10110101",
   "01101000",
   "11111011",
   "00001010",
   "11100100",
   "11110000",
   "00001010",
   "00101100",
   "00011010",
   "11100000",
   "01101000",
   "00011000",
   "00110101",
   "11011101",
   "11110111",
   "11010100",
   "00001010",
   "00101000",
   "00011010",
   "01001100",
   "10110011",
   "11111000",
   "00110001",
   "00011100",
   "00110110",
   "11101110",
   "01010111",
   "11101100",
   "00000001",
   "11111110",
   "01100100",
   "11111000",
   "00101001",
   "00101001",
   "00101110",
   "00010000",
   "11111110",
   "11100110",
   "11001010",
   "00000110",
   "10100001",
   "11000111",
   "00000110",
   "01001110",
   "11010111",
   "00011001",
   "10011000",
   "11111010",
   "00100111",
   "00101000",
   "00000000",
   "01001110",
   "10110111",
   "00010011",
   "00100000",
   "00101110",
   "00000111",
   "00100100",
   "11111100",
   "11110110",
   "11011010",
   "00110011",
   "11011101",
   "01000100",
   "00110000",
   "00000101",
   "11111000",
   "01010100",
   "10100011",
   "00000010",
   "11111001",
   "00000010",
   "00110010",
   "11011010",
   "00010110",
   "11010110",
   "00000010",
   "00111100",
   "01001010",
   "11111010",
   "10100110",
   "11011101",
   "00000010",
   "11100010",
   "00001111",
   "11100101",
   "10111010",
   "11101100",
   "00011101",
   "11110001",
   "10111000",
   "00010000",
   "11010001",
   "11010010",
   "10001110",
   "11000100",
   "11101010",
   "10110010",
   "00000111",
   "11011100",
   "00100110",
   "00001010",
   "01010001",
   "01010000",
   "00111010",
   "00010100",
   "11111001",
   "11111000",
   "00011110",
   "00001000",
   "11011110",
   "11100110",
   "11010101",
   "11000110",
   "00110000",
   "00000110",
   "10110001",
   "01010110",
   "11111011",
   "00011010",
   "11101100",
   "00000111",
   "10100101",
   "11011010",
   "10101001",
   "11011000",
   "01111100",
   "00111100",
   "10110101",
   "11110011",
   "11100100",
   "10001100",
   "11111101",
   "00011111",
   "00000100",
   "00011110",
   "00110110",
   "01001011",
   "00001000",
   "00010110",
   "00101100",
   "11010101",
   "11100001",
   "00000110",
   "00101011",
   "11000000",
   "00000110",
   "11001110",
   "00001100",
   "11111110",
   "00001001",
   "01000110",
   "00110010",
   "11111001",
   "00011101",
   "11101110",
   "00000111",
   "11101010",
   "10010010",
	others => "00000000"
   );
begin
   -- addr register to infer block RAM
   process (clk)
   begin
      if (rising_edge(clk)) then
        addr_reg <= addr;
      end if;
   end process;
   data0 <= signed(ROM(to_integer(unsigned(addr_reg))));
   data1 <= signed(ROM(to_integer(unsigned(addr_reg))+1));
   data2 <= signed(ROM(to_integer(unsigned(addr_reg))+2));
   data3 <= signed(ROM(to_integer(unsigned(addr_reg))+3));
   data4 <= signed(ROM(to_integer(unsigned(addr_reg))+4));
   data5 <= signed(ROM(to_integer(unsigned(addr_reg))+5));
   data6 <= signed(ROM(to_integer(unsigned(addr_reg))+6));
   data7 <= signed(ROM(to_integer(unsigned(addr_reg))+7));

end arc;
